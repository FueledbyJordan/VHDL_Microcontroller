LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MEMORY IS
PORT(
address : IN STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
dataout : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
datain : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
readwrite : IN STD_LOGIC;-- := '0';   --read is 0, write is 1
clk : in STD_LOGIC := '0';
rst : in STD_LOGIC := '0'
);
END ENTITY;

ARCHITECTURE BEV OF MEMORY IS
TYPE MEM_2048 IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL MEMORY : MEM_2048 := (OTHERS => "00000000");
SHARED VARIABLE ADDR : INTEGER RANGE 0 TO 255;
BEGIN
MEMORY(0) <= "00000000";
MEMORY(1) <= "11100100";
MEMORY(2) <= "00000000";
MEMORY(3) <= "11100000";
MEMORY(4) <= "10000000";
MEMORY(5) <= "01001000";
MEMORY(6) <= "10001000";
MEMORY(7) <= "00001110";
MEMORY(8) <= "00100110";
MEMORY(9) <= "11101100";
MEMORY(10) <= "00000001";
MEMORY(11) <= "00100011";
MEMORY(12) <= "11111111";
MEMORY(13) <= "00000101";
MEMORY(14) <= "11010100";
MEMORY(15) <= "01000000";
MEMORY(16) <= "11111111";
MEMORY(17) <= "00010000";
MEMORY(18) <= "00000000";
MEMORY(128) <= "10000000";
MEMORY(129) <= "10000001";
MEMORY(130) <= "10000010";
MEMORY(131) <= "10000011";
MEMORY(132) <= "10000100";
MEMORY(133) <= "10000101";
MEMORY(134) <= "10000110";
MEMORY(135) <= "10000111";
MEMORY(136) <= "10001000";
MEMORY(137) <= "10001001";
MEMORY(138) <= "10001010";
MEMORY(139) <= "10001011";
MEMORY(140) <= "10001100";
MEMORY(141) <= "10001101";
MEMORY(142) <= "10001110";
MEMORY(143) <= "10001111";
MEMORY(144) <= "10010000";
MEMORY(145) <= "10010001";
MEMORY(146) <= "10010010";
MEMORY(147) <= "10010011";
MEMORY(148) <= "10010100";
MEMORY(149) <= "10010101";
MEMORY(150) <= "10010110";
MEMORY(151) <= "10010111";
MEMORY(152) <= "10011000";
MEMORY(153) <= "10011001";
MEMORY(154) <= "10011010";
MEMORY(155) <= "10011011";
MEMORY(156) <= "10011100";
MEMORY(157) <= "10011101";
MEMORY(158) <= "10011110";
MEMORY(159) <= "10011111";
PROCESS(ADDRESS, DATAIN, readwrite, clk, rst)
BEGIN
IF(rising_edge(clk)) THEN
IF(rst='1') THEN
dataout <= "00000000";
ELSE
ADDR:=CONV_INTEGER(ADDRESS);
IF(readwrite='1')THEN
MEMORY(ADDR)<=datain;
ELSE
dataout<=MEMORY(ADDR);
END IF;
END IF;
END IF;
END PROCESS;
END BEV;
